module ethers

fn main() {
	println('Hello World!')
}
