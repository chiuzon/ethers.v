module ethers

import math.big

