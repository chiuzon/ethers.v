module providers

struct JsonProvider {
	pub mut:
		rpc_url string
}

