module utils


pub fn cut_o_x(str string) string {
	return str[2..str.len]
}