module transactions

pub fn sign_tx_with_private_key() {
	// TODO
}